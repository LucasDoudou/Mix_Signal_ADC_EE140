//Verilog HDL for "EECS151T", "Inverter_test" "functional"


module Inverter_test (input x, output y );
assign y = ~x;
endmodule
